// /*###############################################
// #            DEVICE Test Bench MODULE           #
// ################################################*/

// //include "Device.v";

// module DEVICE_tb();
// /*################## REG ##################*/
// reg CLK_tb;
// reg RST_tb;
// reg FRAME_tb;
// reg [3:0] CBE_tb;
// reg IRDY_tb;
// /*################## NET ##################*/
// wire [31: 0] AD_tb;
// wire TRDY_tb;
// wire DEVSEL_tb;




// //Device D1(); // by position

// initial 
// begin: GENERATE_CLK 
//     CLK_tb <= 1;
//     always
//     begin 
//         #1 // f = ??
//         CLK_tb <= ~CLK_tb;
//     end
// end


// initial 
// begin
// /*################ TEST WRITE OPERATION #################*/

// /*################ TEST READ OPERATION #################*/

// end
// endmodule

