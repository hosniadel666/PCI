/*###############################################
#            DEVICE Test Bench MODULE           #
################################################*/

module DEVICE_tb();

endmodule

